//`timescale 1ns / 1ps

module tb_memory_module;

    reg clk;
    reg rst;

    // ------------------------------------------------
    // INPUTS
    // ------------------------------------------------
    // Matrix A Inputs
    reg [7:0] A11, A12, A13, A14;
    reg [7:0] A21, A22, A23, A24;
    reg [7:0] A31, A32, A33, A34;
    reg [7:0] A41, A42, A43, A44;

    // Filter B Inputs
    reg [7:0] B11, B12, B13;
    reg [7:0] B21, B22, B23;
    reg [7:0] B31, B32, B33;

    // ------------------------------------------------
    // OUTPUTS
    // ------------------------------------------------
    wire [7:0] out_A11, out_A12, out_A13, out_A14;
    wire [7:0] out_A21, out_A22, out_A23, out_A24;
    wire [7:0] out_A31, out_A32, out_A33, out_A34;
    wire [7:0] out_A41, out_A42, out_A43, out_A44;

    wire [7:0] out_B11, out_B12, out_B13;
    wire [7:0] out_B21, out_B22, out_B23;
    wire [7:0] out_B31, out_B32, out_B33;

    // ------------------------------------------------
    // MODULE INSTANCE
    // ------------------------------------------------
    memory_module_2 uut (
        .clk(clk), .rst(rst), 
        .A11(A11), .A12(A12), .A13(A13), .A14(A14),
        .A21(A21), .A22(A22), .A23(A23), .A24(A24),
        .A31(A31), .A32(A32), .A33(A33), .A34(A34),
        .A41(A41), .A42(A42), .A43(A43), .A44(A44),
        .B11(B11), .B12(B12), .B13(B13),
        .B21(B21), .B22(B22), .B23(B23),
        .B31(B31), .B32(B32), .B33(B33),
        .out_A11(out_A11), .out_A12(out_A12), .out_A13(out_A13), .out_A14(out_A14),
        .out_A21(out_A21), .out_A22(out_A22), .out_A23(out_A23), .out_A24(out_A24),
        .out_A31(out_A31), .out_A32(out_A32), .out_A33(out_A33), .out_A34(out_A34),
        .out_A41(out_A41), .out_A42(out_A42), .out_A43(out_A43), .out_A44(out_A44),
        .out_B11(out_B11), .out_B12(out_B12), .out_B13(out_B13),
        .out_B21(out_B21), .out_B22(out_B22), .out_B23(out_B23),
        .out_B31(out_B31), .out_B32(out_B32), .out_B33(out_B33)
    );

    // Fast Clock Generation (Period 2ns)
    always #1 clk = ~clk;

    initial begin
        // ???
        clk = 0;
        rst = 0; 

        // ===========================================================
        // [PHASE 1] ?? ??? ?? (?: 1 ~ 25)
        // ===========================================================
        A11=1;  A12=2;  A13=3;  A14=4;
        A21=5;  A22=6;  A23=7;  A24=8;
        A31=9;  A32=10; A33=11; A34=12;
        A41=13; A42=14; A43=15; A44=16;
        
        B11=17; B12=18; B13=19;
        B21=20; B22=21; B23=22;
        B31=23; B32=24; B33=25;

        #10; // Waveform ??: ??? 1~25 ?? ??

        // ===========================================================
        // [PHASE 2] Reset ?? ?? (rst=1 -> ?? 0)
        // ===========================================================
        rst = 1;

        #10; // Waveform ??: ?? ??? 00000000 (0) ?? ??

        // ===========================================================
        // [PHASE 3] ??? ??? ?? (?: 101 ~ 125)
        // Reset ?? ? ?? ????? ???? ??
        // ===========================================================
        rst = 0; // Reset ??

        A11=101; A12=102; A13=103; A14=104;
        A21=105; A22=106; A23=107; A24=108;
        A31=109; A32=110; A33=111; A34=112;
        A41=113; A42=114; A43=115; A44=116;
        
        B11=117; B12=118; B13=119;
        B21=120; B22=121; B23=122;
        B31=123; B32=124; B33=125;

        #10; // Waveform ??: ??? 101~125 ? ????? ??

        $finish;
    end

endmodule