module top_module (
    input clk,
    input rst,

);


endmodule