module top_module (
    input clk,
    input rst,
    input start,
);




endmodule