module controller (
    input clk,
    input rst,

);

// input 정의(원래는 밖에서 받아야하나 이 모듈에서는 미리 내부에 값들을 하드 코딩)


// controller state 정의


// memory에 input 저장


// conv_pe 모듈 instantiation


// output 결과 처리


// conv_sa2x2 모듈 instantiation


// output 결과 처리


// conv_3x3 모듈 instantiation


// output 결과 처리


// display 결과 처리
endmodule