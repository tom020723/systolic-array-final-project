module seven_segment (
    input [3:0] binary_in,
    output reg [6:0] seg_out
);

endmodule